library verilog;
use verilog.vl_types.all;
entity M8_1E_HXILINX_merge_arrays_mcu is
    port(
        O               : out    vl_logic;
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        D4              : in     vl_logic;
        D5              : in     vl_logic;
        D6              : in     vl_logic;
        D7              : in     vl_logic;
        E               : in     vl_logic;
        S0              : in     vl_logic;
        S1              : in     vl_logic;
        S2              : in     vl_logic
    );
end M8_1E_HXILINX_merge_arrays_mcu;
