library verilog;
use verilog.vl_types.all;
entity ee201_GCD_CEN_tb_v is
end ee201_GCD_CEN_tb_v;
